netcdf simple {
dimensions:
	latitude = 3 ;
	longitude = 2 ;
	time = UNLIMITED ; // (5 currently);
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:units = "minutes since 1994-01-01 00:00:00" ;
		time:long_name = "time" ;
	float latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:point_spacing = "even" ;
		latitude:long_name = "latitude" ;
	float longitude(longitude) ;
  		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:point_spacing = "even" ;
		longitude:long_name = "longitude" ;
	float temp(time, latitude, longitude) ;
		temp:standard_name = "surface_temperature" ;
		temp:long_name = "Surface temperature in degrees C" ;
		temp:units = "deg_C" ;
		temp:_FillValue = 2.e+020f ;
		temp:valid_min = -80.f ;
		temp:valid_max = 60.f ;
		temp:comment = "This parameter may be erroneous." ;

// global attributes:
                :Conventions = "CF-1.0" ;
		:institute = "The British Atmospheric Data Centre." ;
		:source = "Model developed in conjunction with IPLSPSC." ;
		:history = "10 Sep 2002 - Created by hand.\n",
			   "18 Mar 2003 - Modified by feet.\n" ;
		:title = "Model output from imaginary model (temperONETER)." ;
		:comment = "Not very useful data." ;
		:references = "A great report somewhere!" ;

data:

 time = 0.5, 1.5, 2.5, 3.5, 4.5 ;

 latitude = 54.2, 54.4, 54.6 ;

 longitude = 2.0, 2.5 ;

 temp =  34.5,  31.2,  23.7,  19.6,  35.8,  29.2,  24.4, 5.6, 7.2, 8.1,
 18.6,  15.2,  13.1, 4.6, 3.7, 8.2, 9.7, 34.2, 26.7, 28.7,
 2.1, 3.4, 5.6, 7.8, 9.0, 10.2, 11.2, 11.6, 11.7, 11.8 ;
}
